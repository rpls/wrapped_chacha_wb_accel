VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_chacha_wb_accel
  CLASS BLOCK ;
  FOREIGN wrapped_chacha_wb_accel ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.850 346.000 30.410 350.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1.100 350.000 2.300 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 92.900 350.000 94.100 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 102.420 350.000 103.620 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 111.260 350.000 112.460 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 120.780 350.000 121.980 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 129.620 350.000 130.820 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 139.140 350.000 140.340 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 147.980 350.000 149.180 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 157.500 350.000 158.700 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 166.340 350.000 167.540 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 175.860 350.000 177.060 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 9.940 350.000 11.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 185.380 350.000 186.580 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 194.220 350.000 195.420 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 203.740 350.000 204.940 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 212.580 350.000 213.780 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 222.100 350.000 223.300 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 230.940 350.000 232.140 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 240.460 350.000 241.660 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 249.300 350.000 250.500 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 258.820 350.000 260.020 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 268.340 350.000 269.540 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 19.460 350.000 20.660 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 277.180 350.000 278.380 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 286.700 350.000 287.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 295.540 350.000 296.740 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 305.060 350.000 306.260 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 313.900 350.000 315.100 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 323.420 350.000 324.620 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 332.260 350.000 333.460 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 341.780 350.000 342.980 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 28.300 350.000 29.500 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 37.820 350.000 39.020 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 46.660 350.000 47.860 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 56.180 350.000 57.380 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 65.020 350.000 66.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 74.540 350.000 75.740 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 83.380 350.000 84.580 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 7.220 350.000 8.420 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 99.020 350.000 100.220 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 108.540 350.000 109.740 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 117.380 350.000 118.580 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 126.900 350.000 128.100 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 135.740 350.000 136.940 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 145.260 350.000 146.460 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 154.100 350.000 155.300 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 163.620 350.000 164.820 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 172.460 350.000 173.660 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 181.980 350.000 183.180 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 16.060 350.000 17.260 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 191.500 350.000 192.700 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 200.340 350.000 201.540 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 209.860 350.000 211.060 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 218.700 350.000 219.900 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 228.220 350.000 229.420 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 237.060 350.000 238.260 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 246.580 350.000 247.780 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 255.420 350.000 256.620 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 264.940 350.000 266.140 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 274.460 350.000 275.660 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 25.580 350.000 26.780 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 283.300 350.000 284.500 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 292.820 350.000 294.020 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 301.660 350.000 302.860 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 311.180 350.000 312.380 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 320.020 350.000 321.220 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 329.540 350.000 330.740 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 338.380 350.000 339.580 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 347.900 350.000 349.100 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 34.420 350.000 35.620 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 43.940 350.000 45.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 52.780 350.000 53.980 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 62.300 350.000 63.500 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 71.140 350.000 72.340 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 80.660 350.000 81.860 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 90.180 350.000 91.380 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 3.820 350.000 5.020 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 96.300 350.000 97.500 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 105.140 350.000 106.340 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 114.660 350.000 115.860 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 123.500 350.000 124.700 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 133.020 350.000 134.220 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 141.860 350.000 143.060 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 151.380 350.000 152.580 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 160.220 350.000 161.420 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 169.740 350.000 170.940 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 179.260 350.000 180.460 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 13.340 350.000 14.540 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 188.100 350.000 189.300 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 197.620 350.000 198.820 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 206.460 350.000 207.660 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 215.980 350.000 217.180 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 224.820 350.000 226.020 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 234.340 350.000 235.540 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 243.180 350.000 244.380 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 252.700 350.000 253.900 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 261.540 350.000 262.740 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 271.060 350.000 272.260 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 22.180 350.000 23.380 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 280.580 350.000 281.780 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 289.420 350.000 290.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 298.940 350.000 300.140 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 307.780 350.000 308.980 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 317.300 350.000 318.500 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 326.140 350.000 327.340 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 335.660 350.000 336.860 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 344.500 350.000 345.700 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 31.700 350.000 32.900 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 40.540 350.000 41.740 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 50.060 350.000 51.260 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 58.900 350.000 60.100 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 68.420 350.000 69.620 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 77.260 350.000 78.460 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 86.780 350.000 87.980 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.780 4.000 2.980 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.540 4.000 7.740 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.980 4.000 13.180 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.250 0.000 2.810 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.530 0.000 57.090 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 0.000 62.610 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 0.000 68.130 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.090 0.000 73.650 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.610 0.000 79.170 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.130 0.000 84.690 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.650 0.000 90.210 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.170 0.000 95.730 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.690 0.000 101.250 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.750 0.000 106.310 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.310 0.000 7.870 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.270 0.000 111.830 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.790 0.000 117.350 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.310 0.000 122.870 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.830 0.000 128.390 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.350 0.000 133.910 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.870 0.000 139.430 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 0.000 144.950 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.910 0.000 150.470 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.970 0.000 155.530 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.490 0.000 161.050 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.830 0.000 13.390 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.010 0.000 166.570 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.530 0.000 172.090 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.870 0.000 24.430 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.390 0.000 29.950 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 0.000 35.470 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 0.000 40.990 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.950 0.000 46.510 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.470 0.000 52.030 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 0.000 177.610 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.790 0.000 232.350 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.310 0.000 237.870 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.830 0.000 243.390 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.350 0.000 248.910 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.410 0.000 253.970 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.930 0.000 259.490 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.450 0.000 265.010 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 0.000 270.530 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.490 0.000 276.050 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.010 0.000 281.570 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.570 0.000 183.130 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.530 0.000 287.090 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 0.000 292.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 0.000 298.130 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 0.000 303.190 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.150 0.000 308.710 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.670 0.000 314.230 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.190 0.000 319.750 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.710 0.000 325.270 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.230 0.000 330.790 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 0.000 336.310 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.090 0.000 188.650 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 0.000 341.830 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.790 0.000 347.350 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.610 0.000 194.170 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.130 0.000 199.690 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.190 0.000 204.750 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.710 0.000 210.270 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 0.000 215.790 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.750 0.000 221.310 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.270 0.000 226.830 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.700 4.000 185.900 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.380 4.000 237.580 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.820 4.000 243.020 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.260 4.000 248.460 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.020 4.000 253.220 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.460 4.000 258.660 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.900 4.000 264.100 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.340 4.000 269.540 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.100 4.000 274.300 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.540 4.000 279.740 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.980 4.000 285.180 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.460 4.000 190.660 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 288.740 4.000 289.940 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.180 4.000 295.380 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.620 4.000 300.820 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.380 4.000 305.580 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.820 4.000 311.020 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.260 4.000 316.460 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.020 4.000 321.220 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.460 4.000 326.660 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 330.900 4.000 332.100 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.660 4.000 336.860 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.900 4.000 196.100 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.100 4.000 342.300 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.540 4.000 347.740 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.340 4.000 201.540 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.100 4.000 206.300 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.540 4.000 211.740 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.980 4.000 217.180 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.740 4.000 221.940 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.180 4.000 227.380 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.620 4.000 232.820 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.450 346.000 35.010 350.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.250 346.000 2.810 350.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.850 346.000 7.410 350.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.250 346.000 25.810 350.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.450 346.000 58.010 350.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.450 346.000 104.010 350.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.050 346.000 108.610 350.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.650 346.000 113.210 350.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.250 346.000 117.810 350.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.850 346.000 122.410 350.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 346.000 127.010 350.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.050 346.000 131.610 350.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.650 346.000 136.210 350.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.250 346.000 140.810 350.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.850 346.000 145.410 350.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.050 346.000 62.610 350.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.450 346.000 150.010 350.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.050 346.000 154.610 350.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.650 346.000 159.210 350.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.250 346.000 163.810 350.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 346.000 168.410 350.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.450 346.000 173.010 350.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.050 346.000 177.610 350.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.650 346.000 182.210 350.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.250 346.000 186.810 350.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.850 346.000 191.410 350.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.650 346.000 67.210 350.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.450 346.000 196.010 350.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.050 346.000 200.610 350.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.250 346.000 71.810 350.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.850 346.000 76.410 350.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.450 346.000 81.010 350.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 346.000 85.610 350.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.650 346.000 90.210 350.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.250 346.000 94.810 350.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 346.000 99.410 350.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.050 346.000 16.610 350.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 346.000 205.210 350.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 346.000 251.210 350.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.250 346.000 255.810 350.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.850 346.000 260.410 350.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.450 346.000 265.010 350.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.050 346.000 269.610 350.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.650 346.000 274.210 350.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.250 346.000 278.810 350.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.850 346.000 283.410 350.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.450 346.000 288.010 350.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 346.000 292.610 350.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 346.000 209.810 350.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.650 346.000 297.210 350.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.250 346.000 301.810 350.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.850 346.000 306.410 350.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.450 346.000 311.010 350.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.050 346.000 315.610 350.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.650 346.000 320.210 350.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.250 346.000 324.810 350.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.850 346.000 329.410 350.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 346.000 334.010 350.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.050 346.000 338.610 350.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.850 346.000 214.410 350.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.650 346.000 343.210 350.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 346.000 347.810 350.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.450 346.000 219.010 350.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.050 346.000 223.610 350.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.650 346.000 228.210 350.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.250 346.000 232.810 350.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.850 346.000 237.410 350.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.450 346.000 242.010 350.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.050 346.000 246.610 350.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.420 4.000 18.620 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.100 4.000 70.300 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.540 4.000 75.740 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 79.980 4.000 81.180 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.740 4.000 85.940 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.180 4.000 91.380 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.620 4.000 96.820 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.060 4.000 102.260 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.820 4.000 107.020 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.260 4.000 112.460 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.700 4.000 117.900 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.180 4.000 23.380 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.460 4.000 122.660 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.900 4.000 128.100 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.340 4.000 133.540 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.100 4.000 138.300 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.540 4.000 143.740 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 147.980 4.000 149.180 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.740 4.000 153.940 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.180 4.000 159.380 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.620 4.000 164.820 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.380 4.000 169.580 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.620 4.000 28.820 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.820 4.000 175.020 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.260 4.000 180.460 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.060 4.000 34.260 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.820 4.000 39.020 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.260 4.000 44.460 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.700 4.000 49.900 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.460 4.000 54.660 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.900 4.000 60.100 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.340 4.000 65.540 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.050 346.000 39.610 350.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 346.000 44.210 350.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.250 346.000 48.810 350.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.850 346.000 53.410 350.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.450 346.000 12.010 350.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.650 346.000 21.210 350.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 345.315 337.365 ;
      LAYER met1 ;
        RECT 2.370 6.500 347.690 338.260 ;
      LAYER met2 ;
        RECT 3.090 345.720 6.570 348.685 ;
        RECT 7.690 345.720 11.170 348.685 ;
        RECT 12.290 345.720 15.770 348.685 ;
        RECT 16.890 345.720 20.370 348.685 ;
        RECT 21.490 345.720 24.970 348.685 ;
        RECT 26.090 345.720 29.570 348.685 ;
        RECT 30.690 345.720 34.170 348.685 ;
        RECT 35.290 345.720 38.770 348.685 ;
        RECT 39.890 345.720 43.370 348.685 ;
        RECT 44.490 345.720 47.970 348.685 ;
        RECT 49.090 345.720 52.570 348.685 ;
        RECT 53.690 345.720 57.170 348.685 ;
        RECT 58.290 345.720 61.770 348.685 ;
        RECT 62.890 345.720 66.370 348.685 ;
        RECT 67.490 345.720 70.970 348.685 ;
        RECT 72.090 345.720 75.570 348.685 ;
        RECT 76.690 345.720 80.170 348.685 ;
        RECT 81.290 345.720 84.770 348.685 ;
        RECT 85.890 345.720 89.370 348.685 ;
        RECT 90.490 345.720 93.970 348.685 ;
        RECT 95.090 345.720 98.570 348.685 ;
        RECT 99.690 345.720 103.170 348.685 ;
        RECT 104.290 345.720 107.770 348.685 ;
        RECT 108.890 345.720 112.370 348.685 ;
        RECT 113.490 345.720 116.970 348.685 ;
        RECT 118.090 345.720 121.570 348.685 ;
        RECT 122.690 345.720 126.170 348.685 ;
        RECT 127.290 345.720 130.770 348.685 ;
        RECT 131.890 345.720 135.370 348.685 ;
        RECT 136.490 345.720 139.970 348.685 ;
        RECT 141.090 345.720 144.570 348.685 ;
        RECT 145.690 345.720 149.170 348.685 ;
        RECT 150.290 345.720 153.770 348.685 ;
        RECT 154.890 345.720 158.370 348.685 ;
        RECT 159.490 345.720 162.970 348.685 ;
        RECT 164.090 345.720 167.570 348.685 ;
        RECT 168.690 345.720 172.170 348.685 ;
        RECT 173.290 345.720 176.770 348.685 ;
        RECT 177.890 345.720 181.370 348.685 ;
        RECT 182.490 345.720 185.970 348.685 ;
        RECT 187.090 345.720 190.570 348.685 ;
        RECT 191.690 345.720 195.170 348.685 ;
        RECT 196.290 345.720 199.770 348.685 ;
        RECT 200.890 345.720 204.370 348.685 ;
        RECT 205.490 345.720 208.970 348.685 ;
        RECT 210.090 345.720 213.570 348.685 ;
        RECT 214.690 345.720 218.170 348.685 ;
        RECT 219.290 345.720 222.770 348.685 ;
        RECT 223.890 345.720 227.370 348.685 ;
        RECT 228.490 345.720 231.970 348.685 ;
        RECT 233.090 345.720 236.570 348.685 ;
        RECT 237.690 345.720 241.170 348.685 ;
        RECT 242.290 345.720 245.770 348.685 ;
        RECT 246.890 345.720 250.370 348.685 ;
        RECT 251.490 345.720 254.970 348.685 ;
        RECT 256.090 345.720 259.570 348.685 ;
        RECT 260.690 345.720 264.170 348.685 ;
        RECT 265.290 345.720 268.770 348.685 ;
        RECT 269.890 345.720 273.370 348.685 ;
        RECT 274.490 345.720 277.970 348.685 ;
        RECT 279.090 345.720 282.570 348.685 ;
        RECT 283.690 345.720 287.170 348.685 ;
        RECT 288.290 345.720 291.770 348.685 ;
        RECT 292.890 345.720 296.370 348.685 ;
        RECT 297.490 345.720 300.970 348.685 ;
        RECT 302.090 345.720 305.570 348.685 ;
        RECT 306.690 345.720 310.170 348.685 ;
        RECT 311.290 345.720 314.770 348.685 ;
        RECT 315.890 345.720 319.370 348.685 ;
        RECT 320.490 345.720 323.970 348.685 ;
        RECT 325.090 345.720 328.570 348.685 ;
        RECT 329.690 345.720 333.170 348.685 ;
        RECT 334.290 345.720 337.770 348.685 ;
        RECT 338.890 345.720 342.370 348.685 ;
        RECT 343.490 345.720 346.970 348.685 ;
        RECT 2.400 4.280 347.660 345.720 ;
        RECT 3.090 2.195 7.030 4.280 ;
        RECT 8.150 2.195 12.550 4.280 ;
        RECT 13.670 2.195 18.070 4.280 ;
        RECT 19.190 2.195 23.590 4.280 ;
        RECT 24.710 2.195 29.110 4.280 ;
        RECT 30.230 2.195 34.630 4.280 ;
        RECT 35.750 2.195 40.150 4.280 ;
        RECT 41.270 2.195 45.670 4.280 ;
        RECT 46.790 2.195 51.190 4.280 ;
        RECT 52.310 2.195 56.250 4.280 ;
        RECT 57.370 2.195 61.770 4.280 ;
        RECT 62.890 2.195 67.290 4.280 ;
        RECT 68.410 2.195 72.810 4.280 ;
        RECT 73.930 2.195 78.330 4.280 ;
        RECT 79.450 2.195 83.850 4.280 ;
        RECT 84.970 2.195 89.370 4.280 ;
        RECT 90.490 2.195 94.890 4.280 ;
        RECT 96.010 2.195 100.410 4.280 ;
        RECT 101.530 2.195 105.470 4.280 ;
        RECT 106.590 2.195 110.990 4.280 ;
        RECT 112.110 2.195 116.510 4.280 ;
        RECT 117.630 2.195 122.030 4.280 ;
        RECT 123.150 2.195 127.550 4.280 ;
        RECT 128.670 2.195 133.070 4.280 ;
        RECT 134.190 2.195 138.590 4.280 ;
        RECT 139.710 2.195 144.110 4.280 ;
        RECT 145.230 2.195 149.630 4.280 ;
        RECT 150.750 2.195 154.690 4.280 ;
        RECT 155.810 2.195 160.210 4.280 ;
        RECT 161.330 2.195 165.730 4.280 ;
        RECT 166.850 2.195 171.250 4.280 ;
        RECT 172.370 2.195 176.770 4.280 ;
        RECT 177.890 2.195 182.290 4.280 ;
        RECT 183.410 2.195 187.810 4.280 ;
        RECT 188.930 2.195 193.330 4.280 ;
        RECT 194.450 2.195 198.850 4.280 ;
        RECT 199.970 2.195 203.910 4.280 ;
        RECT 205.030 2.195 209.430 4.280 ;
        RECT 210.550 2.195 214.950 4.280 ;
        RECT 216.070 2.195 220.470 4.280 ;
        RECT 221.590 2.195 225.990 4.280 ;
        RECT 227.110 2.195 231.510 4.280 ;
        RECT 232.630 2.195 237.030 4.280 ;
        RECT 238.150 2.195 242.550 4.280 ;
        RECT 243.670 2.195 248.070 4.280 ;
        RECT 249.190 2.195 253.130 4.280 ;
        RECT 254.250 2.195 258.650 4.280 ;
        RECT 259.770 2.195 264.170 4.280 ;
        RECT 265.290 2.195 269.690 4.280 ;
        RECT 270.810 2.195 275.210 4.280 ;
        RECT 276.330 2.195 280.730 4.280 ;
        RECT 281.850 2.195 286.250 4.280 ;
        RECT 287.370 2.195 291.770 4.280 ;
        RECT 292.890 2.195 297.290 4.280 ;
        RECT 298.410 2.195 302.350 4.280 ;
        RECT 303.470 2.195 307.870 4.280 ;
        RECT 308.990 2.195 313.390 4.280 ;
        RECT 314.510 2.195 318.910 4.280 ;
        RECT 320.030 2.195 324.430 4.280 ;
        RECT 325.550 2.195 329.950 4.280 ;
        RECT 331.070 2.195 335.470 4.280 ;
        RECT 336.590 2.195 340.990 4.280 ;
        RECT 342.110 2.195 346.510 4.280 ;
        RECT 347.630 2.195 347.660 4.280 ;
      LAYER met3 ;
        RECT 4.000 348.140 345.600 348.665 ;
        RECT 4.400 347.500 345.600 348.140 ;
        RECT 4.400 346.140 346.000 347.500 ;
        RECT 4.000 346.100 346.000 346.140 ;
        RECT 4.000 344.100 345.600 346.100 ;
        RECT 4.000 343.380 346.000 344.100 ;
        RECT 4.000 342.700 345.600 343.380 ;
        RECT 4.400 341.380 345.600 342.700 ;
        RECT 4.400 340.700 346.000 341.380 ;
        RECT 4.000 339.980 346.000 340.700 ;
        RECT 4.000 337.980 345.600 339.980 ;
        RECT 4.000 337.260 346.000 337.980 ;
        RECT 4.400 335.260 345.600 337.260 ;
        RECT 4.000 333.860 346.000 335.260 ;
        RECT 4.000 332.500 345.600 333.860 ;
        RECT 4.400 331.860 345.600 332.500 ;
        RECT 4.400 331.140 346.000 331.860 ;
        RECT 4.400 330.500 345.600 331.140 ;
        RECT 4.000 329.140 345.600 330.500 ;
        RECT 4.000 327.740 346.000 329.140 ;
        RECT 4.000 327.060 345.600 327.740 ;
        RECT 4.400 325.740 345.600 327.060 ;
        RECT 4.400 325.060 346.000 325.740 ;
        RECT 4.000 325.020 346.000 325.060 ;
        RECT 4.000 323.020 345.600 325.020 ;
        RECT 4.000 321.620 346.000 323.020 ;
        RECT 4.400 319.620 345.600 321.620 ;
        RECT 4.000 318.900 346.000 319.620 ;
        RECT 4.000 316.900 345.600 318.900 ;
        RECT 4.000 316.860 346.000 316.900 ;
        RECT 4.400 315.500 346.000 316.860 ;
        RECT 4.400 314.860 345.600 315.500 ;
        RECT 4.000 313.500 345.600 314.860 ;
        RECT 4.000 312.780 346.000 313.500 ;
        RECT 4.000 311.420 345.600 312.780 ;
        RECT 4.400 310.780 345.600 311.420 ;
        RECT 4.400 309.420 346.000 310.780 ;
        RECT 4.000 309.380 346.000 309.420 ;
        RECT 4.000 307.380 345.600 309.380 ;
        RECT 4.000 306.660 346.000 307.380 ;
        RECT 4.000 305.980 345.600 306.660 ;
        RECT 4.400 304.660 345.600 305.980 ;
        RECT 4.400 303.980 346.000 304.660 ;
        RECT 4.000 303.260 346.000 303.980 ;
        RECT 4.000 301.260 345.600 303.260 ;
        RECT 4.000 301.220 346.000 301.260 ;
        RECT 4.400 300.540 346.000 301.220 ;
        RECT 4.400 299.220 345.600 300.540 ;
        RECT 4.000 298.540 345.600 299.220 ;
        RECT 4.000 297.140 346.000 298.540 ;
        RECT 4.000 295.780 345.600 297.140 ;
        RECT 4.400 295.140 345.600 295.780 ;
        RECT 4.400 294.420 346.000 295.140 ;
        RECT 4.400 293.780 345.600 294.420 ;
        RECT 4.000 292.420 345.600 293.780 ;
        RECT 4.000 291.020 346.000 292.420 ;
        RECT 4.000 290.340 345.600 291.020 ;
        RECT 4.400 289.020 345.600 290.340 ;
        RECT 4.400 288.340 346.000 289.020 ;
        RECT 4.000 288.300 346.000 288.340 ;
        RECT 4.000 286.300 345.600 288.300 ;
        RECT 4.000 285.580 346.000 286.300 ;
        RECT 4.400 284.900 346.000 285.580 ;
        RECT 4.400 283.580 345.600 284.900 ;
        RECT 4.000 282.900 345.600 283.580 ;
        RECT 4.000 282.180 346.000 282.900 ;
        RECT 4.000 280.180 345.600 282.180 ;
        RECT 4.000 280.140 346.000 280.180 ;
        RECT 4.400 278.780 346.000 280.140 ;
        RECT 4.400 278.140 345.600 278.780 ;
        RECT 4.000 276.780 345.600 278.140 ;
        RECT 4.000 276.060 346.000 276.780 ;
        RECT 4.000 274.700 345.600 276.060 ;
        RECT 4.400 274.060 345.600 274.700 ;
        RECT 4.400 272.700 346.000 274.060 ;
        RECT 4.000 272.660 346.000 272.700 ;
        RECT 4.000 270.660 345.600 272.660 ;
        RECT 4.000 269.940 346.000 270.660 ;
        RECT 4.400 267.940 345.600 269.940 ;
        RECT 4.000 266.540 346.000 267.940 ;
        RECT 4.000 264.540 345.600 266.540 ;
        RECT 4.000 264.500 346.000 264.540 ;
        RECT 4.400 263.140 346.000 264.500 ;
        RECT 4.400 262.500 345.600 263.140 ;
        RECT 4.000 261.140 345.600 262.500 ;
        RECT 4.000 260.420 346.000 261.140 ;
        RECT 4.000 259.060 345.600 260.420 ;
        RECT 4.400 258.420 345.600 259.060 ;
        RECT 4.400 257.060 346.000 258.420 ;
        RECT 4.000 257.020 346.000 257.060 ;
        RECT 4.000 255.020 345.600 257.020 ;
        RECT 4.000 254.300 346.000 255.020 ;
        RECT 4.000 253.620 345.600 254.300 ;
        RECT 4.400 252.300 345.600 253.620 ;
        RECT 4.400 251.620 346.000 252.300 ;
        RECT 4.000 250.900 346.000 251.620 ;
        RECT 4.000 248.900 345.600 250.900 ;
        RECT 4.000 248.860 346.000 248.900 ;
        RECT 4.400 248.180 346.000 248.860 ;
        RECT 4.400 246.860 345.600 248.180 ;
        RECT 4.000 246.180 345.600 246.860 ;
        RECT 4.000 244.780 346.000 246.180 ;
        RECT 4.000 243.420 345.600 244.780 ;
        RECT 4.400 242.780 345.600 243.420 ;
        RECT 4.400 242.060 346.000 242.780 ;
        RECT 4.400 241.420 345.600 242.060 ;
        RECT 4.000 240.060 345.600 241.420 ;
        RECT 4.000 238.660 346.000 240.060 ;
        RECT 4.000 237.980 345.600 238.660 ;
        RECT 4.400 236.660 345.600 237.980 ;
        RECT 4.400 235.980 346.000 236.660 ;
        RECT 4.000 235.940 346.000 235.980 ;
        RECT 4.000 233.940 345.600 235.940 ;
        RECT 4.000 233.220 346.000 233.940 ;
        RECT 4.400 232.540 346.000 233.220 ;
        RECT 4.400 231.220 345.600 232.540 ;
        RECT 4.000 230.540 345.600 231.220 ;
        RECT 4.000 229.820 346.000 230.540 ;
        RECT 4.000 227.820 345.600 229.820 ;
        RECT 4.000 227.780 346.000 227.820 ;
        RECT 4.400 226.420 346.000 227.780 ;
        RECT 4.400 225.780 345.600 226.420 ;
        RECT 4.000 224.420 345.600 225.780 ;
        RECT 4.000 223.700 346.000 224.420 ;
        RECT 4.000 222.340 345.600 223.700 ;
        RECT 4.400 221.700 345.600 222.340 ;
        RECT 4.400 220.340 346.000 221.700 ;
        RECT 4.000 220.300 346.000 220.340 ;
        RECT 4.000 218.300 345.600 220.300 ;
        RECT 4.000 217.580 346.000 218.300 ;
        RECT 4.400 215.580 345.600 217.580 ;
        RECT 4.000 214.180 346.000 215.580 ;
        RECT 4.000 212.180 345.600 214.180 ;
        RECT 4.000 212.140 346.000 212.180 ;
        RECT 4.400 211.460 346.000 212.140 ;
        RECT 4.400 210.140 345.600 211.460 ;
        RECT 4.000 209.460 345.600 210.140 ;
        RECT 4.000 208.060 346.000 209.460 ;
        RECT 4.000 206.700 345.600 208.060 ;
        RECT 4.400 206.060 345.600 206.700 ;
        RECT 4.400 205.340 346.000 206.060 ;
        RECT 4.400 204.700 345.600 205.340 ;
        RECT 4.000 203.340 345.600 204.700 ;
        RECT 4.000 201.940 346.000 203.340 ;
        RECT 4.400 199.940 345.600 201.940 ;
        RECT 4.000 199.220 346.000 199.940 ;
        RECT 4.000 197.220 345.600 199.220 ;
        RECT 4.000 196.500 346.000 197.220 ;
        RECT 4.400 195.820 346.000 196.500 ;
        RECT 4.400 194.500 345.600 195.820 ;
        RECT 4.000 193.820 345.600 194.500 ;
        RECT 4.000 193.100 346.000 193.820 ;
        RECT 4.000 191.100 345.600 193.100 ;
        RECT 4.000 191.060 346.000 191.100 ;
        RECT 4.400 189.700 346.000 191.060 ;
        RECT 4.400 189.060 345.600 189.700 ;
        RECT 4.000 187.700 345.600 189.060 ;
        RECT 4.000 186.980 346.000 187.700 ;
        RECT 4.000 186.300 345.600 186.980 ;
        RECT 4.400 184.980 345.600 186.300 ;
        RECT 4.400 184.300 346.000 184.980 ;
        RECT 4.000 183.580 346.000 184.300 ;
        RECT 4.000 181.580 345.600 183.580 ;
        RECT 4.000 180.860 346.000 181.580 ;
        RECT 4.400 178.860 345.600 180.860 ;
        RECT 4.000 177.460 346.000 178.860 ;
        RECT 4.000 175.460 345.600 177.460 ;
        RECT 4.000 175.420 346.000 175.460 ;
        RECT 4.400 174.060 346.000 175.420 ;
        RECT 4.400 173.420 345.600 174.060 ;
        RECT 4.000 172.060 345.600 173.420 ;
        RECT 4.000 171.340 346.000 172.060 ;
        RECT 4.000 169.980 345.600 171.340 ;
        RECT 4.400 169.340 345.600 169.980 ;
        RECT 4.400 167.980 346.000 169.340 ;
        RECT 4.000 167.940 346.000 167.980 ;
        RECT 4.000 165.940 345.600 167.940 ;
        RECT 4.000 165.220 346.000 165.940 ;
        RECT 4.400 163.220 345.600 165.220 ;
        RECT 4.000 161.820 346.000 163.220 ;
        RECT 4.000 159.820 345.600 161.820 ;
        RECT 4.000 159.780 346.000 159.820 ;
        RECT 4.400 159.100 346.000 159.780 ;
        RECT 4.400 157.780 345.600 159.100 ;
        RECT 4.000 157.100 345.600 157.780 ;
        RECT 4.000 155.700 346.000 157.100 ;
        RECT 4.000 154.340 345.600 155.700 ;
        RECT 4.400 153.700 345.600 154.340 ;
        RECT 4.400 152.980 346.000 153.700 ;
        RECT 4.400 152.340 345.600 152.980 ;
        RECT 4.000 150.980 345.600 152.340 ;
        RECT 4.000 149.580 346.000 150.980 ;
        RECT 4.400 147.580 345.600 149.580 ;
        RECT 4.000 146.860 346.000 147.580 ;
        RECT 4.000 144.860 345.600 146.860 ;
        RECT 4.000 144.140 346.000 144.860 ;
        RECT 4.400 143.460 346.000 144.140 ;
        RECT 4.400 142.140 345.600 143.460 ;
        RECT 4.000 141.460 345.600 142.140 ;
        RECT 4.000 140.740 346.000 141.460 ;
        RECT 4.000 138.740 345.600 140.740 ;
        RECT 4.000 138.700 346.000 138.740 ;
        RECT 4.400 137.340 346.000 138.700 ;
        RECT 4.400 136.700 345.600 137.340 ;
        RECT 4.000 135.340 345.600 136.700 ;
        RECT 4.000 134.620 346.000 135.340 ;
        RECT 4.000 133.940 345.600 134.620 ;
        RECT 4.400 132.620 345.600 133.940 ;
        RECT 4.400 131.940 346.000 132.620 ;
        RECT 4.000 131.220 346.000 131.940 ;
        RECT 4.000 129.220 345.600 131.220 ;
        RECT 4.000 128.500 346.000 129.220 ;
        RECT 4.400 126.500 345.600 128.500 ;
        RECT 4.000 125.100 346.000 126.500 ;
        RECT 4.000 123.100 345.600 125.100 ;
        RECT 4.000 123.060 346.000 123.100 ;
        RECT 4.400 122.380 346.000 123.060 ;
        RECT 4.400 121.060 345.600 122.380 ;
        RECT 4.000 120.380 345.600 121.060 ;
        RECT 4.000 118.980 346.000 120.380 ;
        RECT 4.000 118.300 345.600 118.980 ;
        RECT 4.400 116.980 345.600 118.300 ;
        RECT 4.400 116.300 346.000 116.980 ;
        RECT 4.000 116.260 346.000 116.300 ;
        RECT 4.000 114.260 345.600 116.260 ;
        RECT 4.000 112.860 346.000 114.260 ;
        RECT 4.400 110.860 345.600 112.860 ;
        RECT 4.000 110.140 346.000 110.860 ;
        RECT 4.000 108.140 345.600 110.140 ;
        RECT 4.000 107.420 346.000 108.140 ;
        RECT 4.400 106.740 346.000 107.420 ;
        RECT 4.400 105.420 345.600 106.740 ;
        RECT 4.000 104.740 345.600 105.420 ;
        RECT 4.000 104.020 346.000 104.740 ;
        RECT 4.000 102.660 345.600 104.020 ;
        RECT 4.400 102.020 345.600 102.660 ;
        RECT 4.400 100.660 346.000 102.020 ;
        RECT 4.000 100.620 346.000 100.660 ;
        RECT 4.000 98.620 345.600 100.620 ;
        RECT 4.000 97.900 346.000 98.620 ;
        RECT 4.000 97.220 345.600 97.900 ;
        RECT 4.400 95.900 345.600 97.220 ;
        RECT 4.400 95.220 346.000 95.900 ;
        RECT 4.000 94.500 346.000 95.220 ;
        RECT 4.000 92.500 345.600 94.500 ;
        RECT 4.000 91.780 346.000 92.500 ;
        RECT 4.400 89.780 345.600 91.780 ;
        RECT 4.000 88.380 346.000 89.780 ;
        RECT 4.000 86.380 345.600 88.380 ;
        RECT 4.000 86.340 346.000 86.380 ;
        RECT 4.400 84.980 346.000 86.340 ;
        RECT 4.400 84.340 345.600 84.980 ;
        RECT 4.000 82.980 345.600 84.340 ;
        RECT 4.000 82.260 346.000 82.980 ;
        RECT 4.000 81.580 345.600 82.260 ;
        RECT 4.400 80.260 345.600 81.580 ;
        RECT 4.400 79.580 346.000 80.260 ;
        RECT 4.000 78.860 346.000 79.580 ;
        RECT 4.000 76.860 345.600 78.860 ;
        RECT 4.000 76.140 346.000 76.860 ;
        RECT 4.400 74.140 345.600 76.140 ;
        RECT 4.000 72.740 346.000 74.140 ;
        RECT 4.000 70.740 345.600 72.740 ;
        RECT 4.000 70.700 346.000 70.740 ;
        RECT 4.400 70.020 346.000 70.700 ;
        RECT 4.400 68.700 345.600 70.020 ;
        RECT 4.000 68.020 345.600 68.700 ;
        RECT 4.000 66.620 346.000 68.020 ;
        RECT 4.000 65.940 345.600 66.620 ;
        RECT 4.400 64.620 345.600 65.940 ;
        RECT 4.400 63.940 346.000 64.620 ;
        RECT 4.000 63.900 346.000 63.940 ;
        RECT 4.000 61.900 345.600 63.900 ;
        RECT 4.000 60.500 346.000 61.900 ;
        RECT 4.400 58.500 345.600 60.500 ;
        RECT 4.000 57.780 346.000 58.500 ;
        RECT 4.000 55.780 345.600 57.780 ;
        RECT 4.000 55.060 346.000 55.780 ;
        RECT 4.400 54.380 346.000 55.060 ;
        RECT 4.400 53.060 345.600 54.380 ;
        RECT 4.000 52.380 345.600 53.060 ;
        RECT 4.000 51.660 346.000 52.380 ;
        RECT 4.000 50.300 345.600 51.660 ;
        RECT 4.400 49.660 345.600 50.300 ;
        RECT 4.400 48.300 346.000 49.660 ;
        RECT 4.000 48.260 346.000 48.300 ;
        RECT 4.000 46.260 345.600 48.260 ;
        RECT 4.000 45.540 346.000 46.260 ;
        RECT 4.000 44.860 345.600 45.540 ;
        RECT 4.400 43.540 345.600 44.860 ;
        RECT 4.400 42.860 346.000 43.540 ;
        RECT 4.000 42.140 346.000 42.860 ;
        RECT 4.000 40.140 345.600 42.140 ;
        RECT 4.000 39.420 346.000 40.140 ;
        RECT 4.400 37.420 345.600 39.420 ;
        RECT 4.000 36.020 346.000 37.420 ;
        RECT 4.000 34.660 345.600 36.020 ;
        RECT 4.400 34.020 345.600 34.660 ;
        RECT 4.400 33.300 346.000 34.020 ;
        RECT 4.400 32.660 345.600 33.300 ;
        RECT 4.000 31.300 345.600 32.660 ;
        RECT 4.000 29.900 346.000 31.300 ;
        RECT 4.000 29.220 345.600 29.900 ;
        RECT 4.400 27.900 345.600 29.220 ;
        RECT 4.400 27.220 346.000 27.900 ;
        RECT 4.000 27.180 346.000 27.220 ;
        RECT 4.000 25.180 345.600 27.180 ;
        RECT 4.000 23.780 346.000 25.180 ;
        RECT 4.400 21.780 345.600 23.780 ;
        RECT 4.000 21.060 346.000 21.780 ;
        RECT 4.000 19.060 345.600 21.060 ;
        RECT 4.000 19.020 346.000 19.060 ;
        RECT 4.400 17.660 346.000 19.020 ;
        RECT 4.400 17.020 345.600 17.660 ;
        RECT 4.000 15.660 345.600 17.020 ;
        RECT 4.000 14.940 346.000 15.660 ;
        RECT 4.000 13.580 345.600 14.940 ;
        RECT 4.400 12.940 345.600 13.580 ;
        RECT 4.400 11.580 346.000 12.940 ;
        RECT 4.000 11.540 346.000 11.580 ;
        RECT 4.000 9.540 345.600 11.540 ;
        RECT 4.000 8.820 346.000 9.540 ;
        RECT 4.000 8.140 345.600 8.820 ;
        RECT 4.400 6.820 345.600 8.140 ;
        RECT 4.400 6.140 346.000 6.820 ;
        RECT 4.000 5.420 346.000 6.140 ;
        RECT 4.000 3.420 345.600 5.420 ;
        RECT 4.000 3.380 346.000 3.420 ;
        RECT 4.400 2.700 346.000 3.380 ;
        RECT 4.400 2.215 345.600 2.700 ;
      LAYER met4 ;
        RECT 95.975 20.575 97.440 283.385 ;
        RECT 99.840 20.575 174.240 283.385 ;
        RECT 176.640 20.575 192.905 283.385 ;
  END
END wrapped_chacha_wb_accel
END LIBRARY


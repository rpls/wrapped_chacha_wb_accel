VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_chacha_wb_accel
  CLASS BLOCK ;
  FOREIGN wrapped_chacha_wb_accel ;
  ORIGIN 0.000 0.000 ;
  SIZE 350.000 BY 350.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 346.000 30.270 350.000 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 1.400 350.000 2.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 93.200 350.000 93.800 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 102.720 350.000 103.320 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 111.560 350.000 112.160 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 121.080 350.000 121.680 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 129.920 350.000 130.520 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 139.440 350.000 140.040 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 148.280 350.000 148.880 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 157.800 350.000 158.400 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 166.640 350.000 167.240 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 176.160 350.000 176.760 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 10.240 350.000 10.840 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 185.680 350.000 186.280 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 194.520 350.000 195.120 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 204.040 350.000 204.640 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 212.880 350.000 213.480 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 222.400 350.000 223.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 231.240 350.000 231.840 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 240.760 350.000 241.360 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 249.600 350.000 250.200 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 259.120 350.000 259.720 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 268.640 350.000 269.240 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 19.760 350.000 20.360 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 277.480 350.000 278.080 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 287.000 350.000 287.600 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 295.840 350.000 296.440 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 305.360 350.000 305.960 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 314.200 350.000 314.800 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 323.720 350.000 324.320 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 332.560 350.000 333.160 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 342.080 350.000 342.680 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 28.600 350.000 29.200 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 38.120 350.000 38.720 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 46.960 350.000 47.560 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 56.480 350.000 57.080 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 65.320 350.000 65.920 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 74.840 350.000 75.440 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 83.680 350.000 84.280 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 7.520 350.000 8.120 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 99.320 350.000 99.920 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 108.840 350.000 109.440 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 117.680 350.000 118.280 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 127.200 350.000 127.800 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 136.040 350.000 136.640 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 145.560 350.000 146.160 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 154.400 350.000 155.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 163.920 350.000 164.520 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 172.760 350.000 173.360 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 182.280 350.000 182.880 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 16.360 350.000 16.960 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 191.800 350.000 192.400 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 200.640 350.000 201.240 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 210.160 350.000 210.760 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 219.000 350.000 219.600 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 228.520 350.000 229.120 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 237.360 350.000 237.960 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 246.880 350.000 247.480 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 255.720 350.000 256.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 265.240 350.000 265.840 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 274.760 350.000 275.360 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 25.880 350.000 26.480 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 283.600 350.000 284.200 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 293.120 350.000 293.720 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 301.960 350.000 302.560 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 311.480 350.000 312.080 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 320.320 350.000 320.920 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 329.840 350.000 330.440 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 338.680 350.000 339.280 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 348.200 350.000 348.800 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 34.720 350.000 35.320 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 44.240 350.000 44.840 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 53.080 350.000 53.680 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 62.600 350.000 63.200 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 71.440 350.000 72.040 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 80.960 350.000 81.560 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 90.480 350.000 91.080 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 4.120 350.000 4.720 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 96.600 350.000 97.200 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 105.440 350.000 106.040 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 114.960 350.000 115.560 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 123.800 350.000 124.400 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 133.320 350.000 133.920 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 142.160 350.000 142.760 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 151.680 350.000 152.280 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 160.520 350.000 161.120 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 170.040 350.000 170.640 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 179.560 350.000 180.160 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 13.640 350.000 14.240 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 188.400 350.000 189.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 197.920 350.000 198.520 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 206.760 350.000 207.360 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 216.280 350.000 216.880 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 225.120 350.000 225.720 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 234.640 350.000 235.240 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 243.480 350.000 244.080 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 253.000 350.000 253.600 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 261.840 350.000 262.440 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 271.360 350.000 271.960 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 22.480 350.000 23.080 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 280.880 350.000 281.480 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 289.720 350.000 290.320 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 299.240 350.000 299.840 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 308.080 350.000 308.680 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 317.600 350.000 318.200 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 326.440 350.000 327.040 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 335.960 350.000 336.560 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 344.800 350.000 345.400 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 32.000 350.000 32.600 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 40.840 350.000 41.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 50.360 350.000 50.960 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 59.200 350.000 59.800 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 68.720 350.000 69.320 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 77.560 350.000 78.160 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 346.000 87.080 350.000 87.680 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 0.000 128.250 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.490 0.000 133.770 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 0.000 150.330 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 0.000 166.430 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 0.000 171.950 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 0.000 248.770 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 0.000 253.830 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.070 0.000 259.350 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 0.000 281.430 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 0.000 182.990 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.710 0.000 297.990 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.810 0.000 314.090 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.330 0.000 319.610 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.370 0.000 330.650 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.890 0.000 336.170 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.930 0.000 347.210 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.000 4.000 185.600 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 236.680 4.000 237.280 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.200 4.000 263.800 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.920 4.000 300.520 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 195.200 4.000 195.800 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END la_oenb[31]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END la_oenb[3]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END la_oenb[5]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 221.040 4.000 221.640 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 226.480 4.000 227.080 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 346.000 34.870 350.000 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 337.520 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 337.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 337.520 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 346.000 2.670 350.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 346.000 7.270 350.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 346.000 25.670 350.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 346.000 57.870 350.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 346.000 103.870 350.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 346.000 108.470 350.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 346.000 113.070 350.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 346.000 117.670 350.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 346.000 122.270 350.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 346.000 126.870 350.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 346.000 131.470 350.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 346.000 136.070 350.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 346.000 140.670 350.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 346.000 145.270 350.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 346.000 62.470 350.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 346.000 149.870 350.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 346.000 154.470 350.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 346.000 159.070 350.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.390 346.000 163.670 350.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 346.000 168.270 350.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 346.000 172.870 350.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 346.000 177.470 350.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 346.000 182.070 350.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 346.000 186.670 350.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 346.000 191.270 350.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.790 346.000 67.070 350.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 195.590 346.000 195.870 350.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 346.000 200.470 350.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 346.000 71.670 350.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 346.000 76.270 350.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 346.000 80.870 350.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 346.000 85.470 350.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 346.000 90.070 350.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 346.000 94.670 350.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 346.000 99.270 350.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 346.000 16.470 350.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 346.000 205.070 350.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 346.000 251.070 350.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.390 346.000 255.670 350.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 346.000 260.270 350.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 346.000 264.870 350.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 346.000 269.470 350.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 346.000 274.070 350.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 346.000 278.670 350.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 346.000 283.270 350.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 346.000 287.870 350.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.190 346.000 292.470 350.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 346.000 209.670 350.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 346.000 297.070 350.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 346.000 301.670 350.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 346.000 306.270 350.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 346.000 310.870 350.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 346.000 315.470 350.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 346.000 320.070 350.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 346.000 324.670 350.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.990 346.000 329.270 350.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 346.000 333.870 350.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 346.000 338.470 350.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.990 346.000 214.270 350.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 346.000 343.070 350.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 346.000 347.670 350.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.590 346.000 218.870 350.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 346.000 223.470 350.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 346.000 228.070 350.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 346.000 232.670 350.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.990 346.000 237.270 350.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 346.000 241.870 350.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 346.000 246.470 350.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 69.400 4.000 70.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.920 4.000 96.520 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 121.760 4.000 122.360 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 346.000 39.470 350.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 346.000 44.070 350.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 346.000 48.670 350.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 346.000 53.270 350.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 346.000 11.870 350.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 346.000 21.070 350.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 345.315 337.365 ;
      LAYER met1 ;
        RECT 2.370 6.500 347.690 338.260 ;
      LAYER met2 ;
        RECT 2.950 345.720 6.710 348.685 ;
        RECT 7.550 345.720 11.310 348.685 ;
        RECT 12.150 345.720 15.910 348.685 ;
        RECT 16.750 345.720 20.510 348.685 ;
        RECT 21.350 345.720 25.110 348.685 ;
        RECT 25.950 345.720 29.710 348.685 ;
        RECT 30.550 345.720 34.310 348.685 ;
        RECT 35.150 345.720 38.910 348.685 ;
        RECT 39.750 345.720 43.510 348.685 ;
        RECT 44.350 345.720 48.110 348.685 ;
        RECT 48.950 345.720 52.710 348.685 ;
        RECT 53.550 345.720 57.310 348.685 ;
        RECT 58.150 345.720 61.910 348.685 ;
        RECT 62.750 345.720 66.510 348.685 ;
        RECT 67.350 345.720 71.110 348.685 ;
        RECT 71.950 345.720 75.710 348.685 ;
        RECT 76.550 345.720 80.310 348.685 ;
        RECT 81.150 345.720 84.910 348.685 ;
        RECT 85.750 345.720 89.510 348.685 ;
        RECT 90.350 345.720 94.110 348.685 ;
        RECT 94.950 345.720 98.710 348.685 ;
        RECT 99.550 345.720 103.310 348.685 ;
        RECT 104.150 345.720 107.910 348.685 ;
        RECT 108.750 345.720 112.510 348.685 ;
        RECT 113.350 345.720 117.110 348.685 ;
        RECT 117.950 345.720 121.710 348.685 ;
        RECT 122.550 345.720 126.310 348.685 ;
        RECT 127.150 345.720 130.910 348.685 ;
        RECT 131.750 345.720 135.510 348.685 ;
        RECT 136.350 345.720 140.110 348.685 ;
        RECT 140.950 345.720 144.710 348.685 ;
        RECT 145.550 345.720 149.310 348.685 ;
        RECT 150.150 345.720 153.910 348.685 ;
        RECT 154.750 345.720 158.510 348.685 ;
        RECT 159.350 345.720 163.110 348.685 ;
        RECT 163.950 345.720 167.710 348.685 ;
        RECT 168.550 345.720 172.310 348.685 ;
        RECT 173.150 345.720 176.910 348.685 ;
        RECT 177.750 345.720 181.510 348.685 ;
        RECT 182.350 345.720 186.110 348.685 ;
        RECT 186.950 345.720 190.710 348.685 ;
        RECT 191.550 345.720 195.310 348.685 ;
        RECT 196.150 345.720 199.910 348.685 ;
        RECT 200.750 345.720 204.510 348.685 ;
        RECT 205.350 345.720 209.110 348.685 ;
        RECT 209.950 345.720 213.710 348.685 ;
        RECT 214.550 345.720 218.310 348.685 ;
        RECT 219.150 345.720 222.910 348.685 ;
        RECT 223.750 345.720 227.510 348.685 ;
        RECT 228.350 345.720 232.110 348.685 ;
        RECT 232.950 345.720 236.710 348.685 ;
        RECT 237.550 345.720 241.310 348.685 ;
        RECT 242.150 345.720 245.910 348.685 ;
        RECT 246.750 345.720 250.510 348.685 ;
        RECT 251.350 345.720 255.110 348.685 ;
        RECT 255.950 345.720 259.710 348.685 ;
        RECT 260.550 345.720 264.310 348.685 ;
        RECT 265.150 345.720 268.910 348.685 ;
        RECT 269.750 345.720 273.510 348.685 ;
        RECT 274.350 345.720 278.110 348.685 ;
        RECT 278.950 345.720 282.710 348.685 ;
        RECT 283.550 345.720 287.310 348.685 ;
        RECT 288.150 345.720 291.910 348.685 ;
        RECT 292.750 345.720 296.510 348.685 ;
        RECT 297.350 345.720 301.110 348.685 ;
        RECT 301.950 345.720 305.710 348.685 ;
        RECT 306.550 345.720 310.310 348.685 ;
        RECT 311.150 345.720 314.910 348.685 ;
        RECT 315.750 345.720 319.510 348.685 ;
        RECT 320.350 345.720 324.110 348.685 ;
        RECT 324.950 345.720 328.710 348.685 ;
        RECT 329.550 345.720 333.310 348.685 ;
        RECT 334.150 345.720 337.910 348.685 ;
        RECT 338.750 345.720 342.510 348.685 ;
        RECT 343.350 345.720 347.110 348.685 ;
        RECT 2.400 4.280 347.660 345.720 ;
        RECT 2.950 2.195 7.170 4.280 ;
        RECT 8.010 2.195 12.690 4.280 ;
        RECT 13.530 2.195 18.210 4.280 ;
        RECT 19.050 2.195 23.730 4.280 ;
        RECT 24.570 2.195 29.250 4.280 ;
        RECT 30.090 2.195 34.770 4.280 ;
        RECT 35.610 2.195 40.290 4.280 ;
        RECT 41.130 2.195 45.810 4.280 ;
        RECT 46.650 2.195 51.330 4.280 ;
        RECT 52.170 2.195 56.390 4.280 ;
        RECT 57.230 2.195 61.910 4.280 ;
        RECT 62.750 2.195 67.430 4.280 ;
        RECT 68.270 2.195 72.950 4.280 ;
        RECT 73.790 2.195 78.470 4.280 ;
        RECT 79.310 2.195 83.990 4.280 ;
        RECT 84.830 2.195 89.510 4.280 ;
        RECT 90.350 2.195 95.030 4.280 ;
        RECT 95.870 2.195 100.550 4.280 ;
        RECT 101.390 2.195 105.610 4.280 ;
        RECT 106.450 2.195 111.130 4.280 ;
        RECT 111.970 2.195 116.650 4.280 ;
        RECT 117.490 2.195 122.170 4.280 ;
        RECT 123.010 2.195 127.690 4.280 ;
        RECT 128.530 2.195 133.210 4.280 ;
        RECT 134.050 2.195 138.730 4.280 ;
        RECT 139.570 2.195 144.250 4.280 ;
        RECT 145.090 2.195 149.770 4.280 ;
        RECT 150.610 2.195 154.830 4.280 ;
        RECT 155.670 2.195 160.350 4.280 ;
        RECT 161.190 2.195 165.870 4.280 ;
        RECT 166.710 2.195 171.390 4.280 ;
        RECT 172.230 2.195 176.910 4.280 ;
        RECT 177.750 2.195 182.430 4.280 ;
        RECT 183.270 2.195 187.950 4.280 ;
        RECT 188.790 2.195 193.470 4.280 ;
        RECT 194.310 2.195 198.990 4.280 ;
        RECT 199.830 2.195 204.050 4.280 ;
        RECT 204.890 2.195 209.570 4.280 ;
        RECT 210.410 2.195 215.090 4.280 ;
        RECT 215.930 2.195 220.610 4.280 ;
        RECT 221.450 2.195 226.130 4.280 ;
        RECT 226.970 2.195 231.650 4.280 ;
        RECT 232.490 2.195 237.170 4.280 ;
        RECT 238.010 2.195 242.690 4.280 ;
        RECT 243.530 2.195 248.210 4.280 ;
        RECT 249.050 2.195 253.270 4.280 ;
        RECT 254.110 2.195 258.790 4.280 ;
        RECT 259.630 2.195 264.310 4.280 ;
        RECT 265.150 2.195 269.830 4.280 ;
        RECT 270.670 2.195 275.350 4.280 ;
        RECT 276.190 2.195 280.870 4.280 ;
        RECT 281.710 2.195 286.390 4.280 ;
        RECT 287.230 2.195 291.910 4.280 ;
        RECT 292.750 2.195 297.430 4.280 ;
        RECT 298.270 2.195 302.490 4.280 ;
        RECT 303.330 2.195 308.010 4.280 ;
        RECT 308.850 2.195 313.530 4.280 ;
        RECT 314.370 2.195 319.050 4.280 ;
        RECT 319.890 2.195 324.570 4.280 ;
        RECT 325.410 2.195 330.090 4.280 ;
        RECT 330.930 2.195 335.610 4.280 ;
        RECT 336.450 2.195 341.130 4.280 ;
        RECT 341.970 2.195 346.650 4.280 ;
        RECT 347.490 2.195 347.660 4.280 ;
      LAYER met3 ;
        RECT 4.000 347.840 345.600 348.665 ;
        RECT 4.400 347.800 345.600 347.840 ;
        RECT 4.400 346.440 346.000 347.800 ;
        RECT 4.000 345.800 346.000 346.440 ;
        RECT 4.000 344.400 345.600 345.800 ;
        RECT 4.000 343.080 346.000 344.400 ;
        RECT 4.000 342.400 345.600 343.080 ;
        RECT 4.400 341.680 345.600 342.400 ;
        RECT 4.400 341.000 346.000 341.680 ;
        RECT 4.000 339.680 346.000 341.000 ;
        RECT 4.000 338.280 345.600 339.680 ;
        RECT 4.000 336.960 346.000 338.280 ;
        RECT 4.400 335.560 345.600 336.960 ;
        RECT 4.000 333.560 346.000 335.560 ;
        RECT 4.000 332.200 345.600 333.560 ;
        RECT 4.400 332.160 345.600 332.200 ;
        RECT 4.400 330.840 346.000 332.160 ;
        RECT 4.400 330.800 345.600 330.840 ;
        RECT 4.000 329.440 345.600 330.800 ;
        RECT 4.000 327.440 346.000 329.440 ;
        RECT 4.000 326.760 345.600 327.440 ;
        RECT 4.400 326.040 345.600 326.760 ;
        RECT 4.400 325.360 346.000 326.040 ;
        RECT 4.000 324.720 346.000 325.360 ;
        RECT 4.000 323.320 345.600 324.720 ;
        RECT 4.000 321.320 346.000 323.320 ;
        RECT 4.400 319.920 345.600 321.320 ;
        RECT 4.000 318.600 346.000 319.920 ;
        RECT 4.000 317.200 345.600 318.600 ;
        RECT 4.000 316.560 346.000 317.200 ;
        RECT 4.400 315.200 346.000 316.560 ;
        RECT 4.400 315.160 345.600 315.200 ;
        RECT 4.000 313.800 345.600 315.160 ;
        RECT 4.000 312.480 346.000 313.800 ;
        RECT 4.000 311.120 345.600 312.480 ;
        RECT 4.400 311.080 345.600 311.120 ;
        RECT 4.400 309.720 346.000 311.080 ;
        RECT 4.000 309.080 346.000 309.720 ;
        RECT 4.000 307.680 345.600 309.080 ;
        RECT 4.000 306.360 346.000 307.680 ;
        RECT 4.000 305.680 345.600 306.360 ;
        RECT 4.400 304.960 345.600 305.680 ;
        RECT 4.400 304.280 346.000 304.960 ;
        RECT 4.000 302.960 346.000 304.280 ;
        RECT 4.000 301.560 345.600 302.960 ;
        RECT 4.000 300.920 346.000 301.560 ;
        RECT 4.400 300.240 346.000 300.920 ;
        RECT 4.400 299.520 345.600 300.240 ;
        RECT 4.000 298.840 345.600 299.520 ;
        RECT 4.000 296.840 346.000 298.840 ;
        RECT 4.000 295.480 345.600 296.840 ;
        RECT 4.400 295.440 345.600 295.480 ;
        RECT 4.400 294.120 346.000 295.440 ;
        RECT 4.400 294.080 345.600 294.120 ;
        RECT 4.000 292.720 345.600 294.080 ;
        RECT 4.000 290.720 346.000 292.720 ;
        RECT 4.000 290.040 345.600 290.720 ;
        RECT 4.400 289.320 345.600 290.040 ;
        RECT 4.400 288.640 346.000 289.320 ;
        RECT 4.000 288.000 346.000 288.640 ;
        RECT 4.000 286.600 345.600 288.000 ;
        RECT 4.000 285.280 346.000 286.600 ;
        RECT 4.400 284.600 346.000 285.280 ;
        RECT 4.400 283.880 345.600 284.600 ;
        RECT 4.000 283.200 345.600 283.880 ;
        RECT 4.000 281.880 346.000 283.200 ;
        RECT 4.000 280.480 345.600 281.880 ;
        RECT 4.000 279.840 346.000 280.480 ;
        RECT 4.400 278.480 346.000 279.840 ;
        RECT 4.400 278.440 345.600 278.480 ;
        RECT 4.000 277.080 345.600 278.440 ;
        RECT 4.000 275.760 346.000 277.080 ;
        RECT 4.000 274.400 345.600 275.760 ;
        RECT 4.400 274.360 345.600 274.400 ;
        RECT 4.400 273.000 346.000 274.360 ;
        RECT 4.000 272.360 346.000 273.000 ;
        RECT 4.000 270.960 345.600 272.360 ;
        RECT 4.000 269.640 346.000 270.960 ;
        RECT 4.400 268.240 345.600 269.640 ;
        RECT 4.000 266.240 346.000 268.240 ;
        RECT 4.000 264.840 345.600 266.240 ;
        RECT 4.000 264.200 346.000 264.840 ;
        RECT 4.400 262.840 346.000 264.200 ;
        RECT 4.400 262.800 345.600 262.840 ;
        RECT 4.000 261.440 345.600 262.800 ;
        RECT 4.000 260.120 346.000 261.440 ;
        RECT 4.000 258.760 345.600 260.120 ;
        RECT 4.400 258.720 345.600 258.760 ;
        RECT 4.400 257.360 346.000 258.720 ;
        RECT 4.000 256.720 346.000 257.360 ;
        RECT 4.000 255.320 345.600 256.720 ;
        RECT 4.000 254.000 346.000 255.320 ;
        RECT 4.000 253.320 345.600 254.000 ;
        RECT 4.400 252.600 345.600 253.320 ;
        RECT 4.400 251.920 346.000 252.600 ;
        RECT 4.000 250.600 346.000 251.920 ;
        RECT 4.000 249.200 345.600 250.600 ;
        RECT 4.000 248.560 346.000 249.200 ;
        RECT 4.400 247.880 346.000 248.560 ;
        RECT 4.400 247.160 345.600 247.880 ;
        RECT 4.000 246.480 345.600 247.160 ;
        RECT 4.000 244.480 346.000 246.480 ;
        RECT 4.000 243.120 345.600 244.480 ;
        RECT 4.400 243.080 345.600 243.120 ;
        RECT 4.400 241.760 346.000 243.080 ;
        RECT 4.400 241.720 345.600 241.760 ;
        RECT 4.000 240.360 345.600 241.720 ;
        RECT 4.000 238.360 346.000 240.360 ;
        RECT 4.000 237.680 345.600 238.360 ;
        RECT 4.400 236.960 345.600 237.680 ;
        RECT 4.400 236.280 346.000 236.960 ;
        RECT 4.000 235.640 346.000 236.280 ;
        RECT 4.000 234.240 345.600 235.640 ;
        RECT 4.000 232.920 346.000 234.240 ;
        RECT 4.400 232.240 346.000 232.920 ;
        RECT 4.400 231.520 345.600 232.240 ;
        RECT 4.000 230.840 345.600 231.520 ;
        RECT 4.000 229.520 346.000 230.840 ;
        RECT 4.000 228.120 345.600 229.520 ;
        RECT 4.000 227.480 346.000 228.120 ;
        RECT 4.400 226.120 346.000 227.480 ;
        RECT 4.400 226.080 345.600 226.120 ;
        RECT 4.000 224.720 345.600 226.080 ;
        RECT 4.000 223.400 346.000 224.720 ;
        RECT 4.000 222.040 345.600 223.400 ;
        RECT 4.400 222.000 345.600 222.040 ;
        RECT 4.400 220.640 346.000 222.000 ;
        RECT 4.000 220.000 346.000 220.640 ;
        RECT 4.000 218.600 345.600 220.000 ;
        RECT 4.000 217.280 346.000 218.600 ;
        RECT 4.400 215.880 345.600 217.280 ;
        RECT 4.000 213.880 346.000 215.880 ;
        RECT 4.000 212.480 345.600 213.880 ;
        RECT 4.000 211.840 346.000 212.480 ;
        RECT 4.400 211.160 346.000 211.840 ;
        RECT 4.400 210.440 345.600 211.160 ;
        RECT 4.000 209.760 345.600 210.440 ;
        RECT 4.000 207.760 346.000 209.760 ;
        RECT 4.000 206.400 345.600 207.760 ;
        RECT 4.400 206.360 345.600 206.400 ;
        RECT 4.400 205.040 346.000 206.360 ;
        RECT 4.400 205.000 345.600 205.040 ;
        RECT 4.000 203.640 345.600 205.000 ;
        RECT 4.000 201.640 346.000 203.640 ;
        RECT 4.400 200.240 345.600 201.640 ;
        RECT 4.000 198.920 346.000 200.240 ;
        RECT 4.000 197.520 345.600 198.920 ;
        RECT 4.000 196.200 346.000 197.520 ;
        RECT 4.400 195.520 346.000 196.200 ;
        RECT 4.400 194.800 345.600 195.520 ;
        RECT 4.000 194.120 345.600 194.800 ;
        RECT 4.000 192.800 346.000 194.120 ;
        RECT 4.000 191.400 345.600 192.800 ;
        RECT 4.000 190.760 346.000 191.400 ;
        RECT 4.400 189.400 346.000 190.760 ;
        RECT 4.400 189.360 345.600 189.400 ;
        RECT 4.000 188.000 345.600 189.360 ;
        RECT 4.000 186.680 346.000 188.000 ;
        RECT 4.000 186.000 345.600 186.680 ;
        RECT 4.400 185.280 345.600 186.000 ;
        RECT 4.400 184.600 346.000 185.280 ;
        RECT 4.000 183.280 346.000 184.600 ;
        RECT 4.000 181.880 345.600 183.280 ;
        RECT 4.000 180.560 346.000 181.880 ;
        RECT 4.400 179.160 345.600 180.560 ;
        RECT 4.000 177.160 346.000 179.160 ;
        RECT 4.000 175.760 345.600 177.160 ;
        RECT 4.000 175.120 346.000 175.760 ;
        RECT 4.400 173.760 346.000 175.120 ;
        RECT 4.400 173.720 345.600 173.760 ;
        RECT 4.000 172.360 345.600 173.720 ;
        RECT 4.000 171.040 346.000 172.360 ;
        RECT 4.000 169.680 345.600 171.040 ;
        RECT 4.400 169.640 345.600 169.680 ;
        RECT 4.400 168.280 346.000 169.640 ;
        RECT 4.000 167.640 346.000 168.280 ;
        RECT 4.000 166.240 345.600 167.640 ;
        RECT 4.000 164.920 346.000 166.240 ;
        RECT 4.400 163.520 345.600 164.920 ;
        RECT 4.000 161.520 346.000 163.520 ;
        RECT 4.000 160.120 345.600 161.520 ;
        RECT 4.000 159.480 346.000 160.120 ;
        RECT 4.400 158.800 346.000 159.480 ;
        RECT 4.400 158.080 345.600 158.800 ;
        RECT 4.000 157.400 345.600 158.080 ;
        RECT 4.000 155.400 346.000 157.400 ;
        RECT 4.000 154.040 345.600 155.400 ;
        RECT 4.400 154.000 345.600 154.040 ;
        RECT 4.400 152.680 346.000 154.000 ;
        RECT 4.400 152.640 345.600 152.680 ;
        RECT 4.000 151.280 345.600 152.640 ;
        RECT 4.000 149.280 346.000 151.280 ;
        RECT 4.400 147.880 345.600 149.280 ;
        RECT 4.000 146.560 346.000 147.880 ;
        RECT 4.000 145.160 345.600 146.560 ;
        RECT 4.000 143.840 346.000 145.160 ;
        RECT 4.400 143.160 346.000 143.840 ;
        RECT 4.400 142.440 345.600 143.160 ;
        RECT 4.000 141.760 345.600 142.440 ;
        RECT 4.000 140.440 346.000 141.760 ;
        RECT 4.000 139.040 345.600 140.440 ;
        RECT 4.000 138.400 346.000 139.040 ;
        RECT 4.400 137.040 346.000 138.400 ;
        RECT 4.400 137.000 345.600 137.040 ;
        RECT 4.000 135.640 345.600 137.000 ;
        RECT 4.000 134.320 346.000 135.640 ;
        RECT 4.000 133.640 345.600 134.320 ;
        RECT 4.400 132.920 345.600 133.640 ;
        RECT 4.400 132.240 346.000 132.920 ;
        RECT 4.000 130.920 346.000 132.240 ;
        RECT 4.000 129.520 345.600 130.920 ;
        RECT 4.000 128.200 346.000 129.520 ;
        RECT 4.400 126.800 345.600 128.200 ;
        RECT 4.000 124.800 346.000 126.800 ;
        RECT 4.000 123.400 345.600 124.800 ;
        RECT 4.000 122.760 346.000 123.400 ;
        RECT 4.400 122.080 346.000 122.760 ;
        RECT 4.400 121.360 345.600 122.080 ;
        RECT 4.000 120.680 345.600 121.360 ;
        RECT 4.000 118.680 346.000 120.680 ;
        RECT 4.000 118.000 345.600 118.680 ;
        RECT 4.400 117.280 345.600 118.000 ;
        RECT 4.400 116.600 346.000 117.280 ;
        RECT 4.000 115.960 346.000 116.600 ;
        RECT 4.000 114.560 345.600 115.960 ;
        RECT 4.000 112.560 346.000 114.560 ;
        RECT 4.400 111.160 345.600 112.560 ;
        RECT 4.000 109.840 346.000 111.160 ;
        RECT 4.000 108.440 345.600 109.840 ;
        RECT 4.000 107.120 346.000 108.440 ;
        RECT 4.400 106.440 346.000 107.120 ;
        RECT 4.400 105.720 345.600 106.440 ;
        RECT 4.000 105.040 345.600 105.720 ;
        RECT 4.000 103.720 346.000 105.040 ;
        RECT 4.000 102.360 345.600 103.720 ;
        RECT 4.400 102.320 345.600 102.360 ;
        RECT 4.400 100.960 346.000 102.320 ;
        RECT 4.000 100.320 346.000 100.960 ;
        RECT 4.000 98.920 345.600 100.320 ;
        RECT 4.000 97.600 346.000 98.920 ;
        RECT 4.000 96.920 345.600 97.600 ;
        RECT 4.400 96.200 345.600 96.920 ;
        RECT 4.400 95.520 346.000 96.200 ;
        RECT 4.000 94.200 346.000 95.520 ;
        RECT 4.000 92.800 345.600 94.200 ;
        RECT 4.000 91.480 346.000 92.800 ;
        RECT 4.400 90.080 345.600 91.480 ;
        RECT 4.000 88.080 346.000 90.080 ;
        RECT 4.000 86.680 345.600 88.080 ;
        RECT 4.000 86.040 346.000 86.680 ;
        RECT 4.400 84.680 346.000 86.040 ;
        RECT 4.400 84.640 345.600 84.680 ;
        RECT 4.000 83.280 345.600 84.640 ;
        RECT 4.000 81.960 346.000 83.280 ;
        RECT 4.000 81.280 345.600 81.960 ;
        RECT 4.400 80.560 345.600 81.280 ;
        RECT 4.400 79.880 346.000 80.560 ;
        RECT 4.000 78.560 346.000 79.880 ;
        RECT 4.000 77.160 345.600 78.560 ;
        RECT 4.000 75.840 346.000 77.160 ;
        RECT 4.400 74.440 345.600 75.840 ;
        RECT 4.000 72.440 346.000 74.440 ;
        RECT 4.000 71.040 345.600 72.440 ;
        RECT 4.000 70.400 346.000 71.040 ;
        RECT 4.400 69.720 346.000 70.400 ;
        RECT 4.400 69.000 345.600 69.720 ;
        RECT 4.000 68.320 345.600 69.000 ;
        RECT 4.000 66.320 346.000 68.320 ;
        RECT 4.000 65.640 345.600 66.320 ;
        RECT 4.400 64.920 345.600 65.640 ;
        RECT 4.400 64.240 346.000 64.920 ;
        RECT 4.000 63.600 346.000 64.240 ;
        RECT 4.000 62.200 345.600 63.600 ;
        RECT 4.000 60.200 346.000 62.200 ;
        RECT 4.400 58.800 345.600 60.200 ;
        RECT 4.000 57.480 346.000 58.800 ;
        RECT 4.000 56.080 345.600 57.480 ;
        RECT 4.000 54.760 346.000 56.080 ;
        RECT 4.400 54.080 346.000 54.760 ;
        RECT 4.400 53.360 345.600 54.080 ;
        RECT 4.000 52.680 345.600 53.360 ;
        RECT 4.000 51.360 346.000 52.680 ;
        RECT 4.000 50.000 345.600 51.360 ;
        RECT 4.400 49.960 345.600 50.000 ;
        RECT 4.400 48.600 346.000 49.960 ;
        RECT 4.000 47.960 346.000 48.600 ;
        RECT 4.000 46.560 345.600 47.960 ;
        RECT 4.000 45.240 346.000 46.560 ;
        RECT 4.000 44.560 345.600 45.240 ;
        RECT 4.400 43.840 345.600 44.560 ;
        RECT 4.400 43.160 346.000 43.840 ;
        RECT 4.000 41.840 346.000 43.160 ;
        RECT 4.000 40.440 345.600 41.840 ;
        RECT 4.000 39.120 346.000 40.440 ;
        RECT 4.400 37.720 345.600 39.120 ;
        RECT 4.000 35.720 346.000 37.720 ;
        RECT 4.000 34.360 345.600 35.720 ;
        RECT 4.400 34.320 345.600 34.360 ;
        RECT 4.400 33.000 346.000 34.320 ;
        RECT 4.400 32.960 345.600 33.000 ;
        RECT 4.000 31.600 345.600 32.960 ;
        RECT 4.000 29.600 346.000 31.600 ;
        RECT 4.000 28.920 345.600 29.600 ;
        RECT 4.400 28.200 345.600 28.920 ;
        RECT 4.400 27.520 346.000 28.200 ;
        RECT 4.000 26.880 346.000 27.520 ;
        RECT 4.000 25.480 345.600 26.880 ;
        RECT 4.000 23.480 346.000 25.480 ;
        RECT 4.400 22.080 345.600 23.480 ;
        RECT 4.000 20.760 346.000 22.080 ;
        RECT 4.000 19.360 345.600 20.760 ;
        RECT 4.000 18.720 346.000 19.360 ;
        RECT 4.400 17.360 346.000 18.720 ;
        RECT 4.400 17.320 345.600 17.360 ;
        RECT 4.000 15.960 345.600 17.320 ;
        RECT 4.000 14.640 346.000 15.960 ;
        RECT 4.000 13.280 345.600 14.640 ;
        RECT 4.400 13.240 345.600 13.280 ;
        RECT 4.400 11.880 346.000 13.240 ;
        RECT 4.000 11.240 346.000 11.880 ;
        RECT 4.000 9.840 345.600 11.240 ;
        RECT 4.000 8.520 346.000 9.840 ;
        RECT 4.000 7.840 345.600 8.520 ;
        RECT 4.400 7.120 345.600 7.840 ;
        RECT 4.400 6.440 346.000 7.120 ;
        RECT 4.000 5.120 346.000 6.440 ;
        RECT 4.000 3.720 345.600 5.120 ;
        RECT 4.000 3.080 346.000 3.720 ;
        RECT 4.400 2.400 346.000 3.080 ;
        RECT 4.400 2.215 345.600 2.400 ;
      LAYER met4 ;
        RECT 95.975 46.415 97.440 283.385 ;
        RECT 99.840 46.415 174.240 283.385 ;
        RECT 176.640 46.415 251.040 283.385 ;
        RECT 253.440 46.415 254.545 283.385 ;
  END
END wrapped_chacha_wb_accel
END LIBRARY

